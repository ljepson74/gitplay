module junk;

   initial begin
      $display(" Atif is a nice boy");
   end

endmodule